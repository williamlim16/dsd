`timescale 1ns / 1ps
`include "Parameter.v"
// fpga4student.com 
// FPGA projects, VHDL projects, Verilog projects 
// Verilog code for RISC Processor 
// Verilog code for data Memory
module Data_Memory(
 input clk,
 // address input, shared by read and write port
 input [15:0]   mem_access_addr,
 
 // write port
 input [15:0]   mem_write_data,
 input     mem_write_en,
 input mem_read,
 // read port
 output [15:0]   mem_read_data
);

reg [`col - 1:0] memory [`row_d - 1:0];
integer f;
wire [2:0] ram_addr=mem_access_addr[2:0];

initial
 begin
	memory[0] = 16'b0000000000000110;
   memory[1] = 16'b0000000000000001;
	memory[2] = 16'b0000000000000001;
	memory[3] = 16'b0000000000000010;
	memory[4] = 16'b0000000000000001;
	memory[5] = 16'b0000000000000010;
	memory[6] = 16'b0000000000000011;
	memory[7] = 16'b0000000000000101;
  `simulation_time;
  
 end

 
 always @(posedge clk) begin
  if (mem_write_en)
   memory[ram_addr] <= mem_write_data;
 end
 assign mem_read_data = (mem_read==1'b1) ? memory[ram_addr]: 16'd0; 

endmodule